// $Id: $
// File name:   mul14.sv
// Created:     4/4/2017
// Author:      Caleb Withers
// Lab Section: 337-02
// Version:     1.0  Initial Design Entry
// Description: Multiply 14

module mul14(
	input wire [7:0]mul14_in,
	output reg [7:0]mul14_out
);

always_comb begin : mul_case
	mul14_out=8'h00;

	case(mul14_in)
		8'h00: mul14_out=8'h00;
		8'h01: mul14_out=8'h0e;
		8'h02: mul14_out=8'h1c;
		8'h03: mul14_out=8'h12;
		8'h04: mul14_out=8'h38;
		8'h05: mul14_out=8'h36;
		8'h06: mul14_out=8'h24;
		8'h07: mul14_out=8'h2a;
		8'h08: mul14_out=8'h70;
		8'h09: mul14_out=8'h7e;
		8'h0a: mul14_out=8'h6c;
		8'h0b: mul14_out=8'h62;
		8'h0c: mul14_out=8'h48;
		8'h0d: mul14_out=8'h46;
		8'h0e: mul14_out=8'h54;
		8'h0f: mul14_out=8'h5a;
		8'h10: mul14_out=8'he0;
		8'h11: mul14_out=8'hee;
		8'h12: mul14_out=8'hfc;
		8'h13: mul14_out=8'hf2;
		8'h14: mul14_out=8'hd8;
		8'h15: mul14_out=8'hd6;
		8'h16: mul14_out=8'hc4;
		8'h17: mul14_out=8'hca;
		8'h18: mul14_out=8'h90;
		8'h19: mul14_out=8'h9e;
		8'h1a: mul14_out=8'h8c;
		8'h1b: mul14_out=8'h82;
		8'h1c: mul14_out=8'ha8;
		8'h1d: mul14_out=8'ha6;
		8'h1e: mul14_out=8'hb4;
		8'h1f: mul14_out=8'hba;
		8'h20: mul14_out=8'hdb;
		8'h21: mul14_out=8'hd5;
		8'h22: mul14_out=8'hc7;
		8'h23: mul14_out=8'hc9;
		8'h24: mul14_out=8'he3;
		8'h25: mul14_out=8'hed;
		8'h26: mul14_out=8'hff;
		8'h27: mul14_out=8'hf1;
		8'h28: mul14_out=8'hab;
		8'h29: mul14_out=8'ha5;
		8'h2a: mul14_out=8'hb7;
		8'h2b: mul14_out=8'hb9;
		8'h2c: mul14_out=8'h93;
		8'h2d: mul14_out=8'h9d;
		8'h2e: mul14_out=8'h8f;
		8'h2f: mul14_out=8'h81;
		8'h30: mul14_out=8'h3b;
		8'h31: mul14_out=8'h35;
		8'h32: mul14_out=8'h27;
		8'h33: mul14_out=8'h29;
		8'h34: mul14_out=8'h03;
		8'h35: mul14_out=8'h0d;
		8'h36: mul14_out=8'h1f;
		8'h37: mul14_out=8'h11;
		8'h38: mul14_out=8'h4b;
		8'h39: mul14_out=8'h45;
		8'h3a: mul14_out=8'h57;
		8'h3b: mul14_out=8'h59;
		8'h3c: mul14_out=8'h73;
		8'h3d: mul14_out=8'h7d;
		8'h3e: mul14_out=8'h6f;
		8'h3f: mul14_out=8'h61;
		8'h40: mul14_out=8'had;
		8'h41: mul14_out=8'ha3;
		8'h42: mul14_out=8'hb1;
		8'h43: mul14_out=8'hbf;
		8'h44: mul14_out=8'h95;
		8'h45: mul14_out=8'h9b;
		8'h46: mul14_out=8'h89;
		8'h47: mul14_out=8'h87;
		8'h48: mul14_out=8'hdd;
		8'h49: mul14_out=8'hd3;
		8'h4a: mul14_out=8'hc1;
		8'h4b: mul14_out=8'hcf;
		8'h4c: mul14_out=8'he5;
		8'h4d: mul14_out=8'heb;
		8'h4e: mul14_out=8'hf9;
		8'h4f: mul14_out=8'hf7;
		8'h50: mul14_out=8'h4d;
		8'h51: mul14_out=8'h43;
		8'h52: mul14_out=8'h51;
		8'h53: mul14_out=8'h5f;
		8'h54: mul14_out=8'h75;
		8'h55: mul14_out=8'h7b;
		8'h56: mul14_out=8'h69;
		8'h57: mul14_out=8'h67;
		8'h58: mul14_out=8'h3d;
		8'h59: mul14_out=8'h33;
		8'h5a: mul14_out=8'h21;
		8'h5b: mul14_out=8'h2f;
		8'h5c: mul14_out=8'h05;
		8'h5d: mul14_out=8'h0b;
		8'h5e: mul14_out=8'h19;
		8'h5f: mul14_out=8'h17;
		8'h60: mul14_out=8'h76;
		8'h61: mul14_out=8'h78;
		8'h62: mul14_out=8'h6a;
		8'h63: mul14_out=8'h64;
		8'h64: mul14_out=8'h4e;
		8'h65: mul14_out=8'h40;
		8'h66: mul14_out=8'h52;
		8'h67: mul14_out=8'h5c;
		8'h68: mul14_out=8'h06;
		8'h69: mul14_out=8'h08;
		8'h6a: mul14_out=8'h1a;
		8'h6b: mul14_out=8'h14;
		8'h6c: mul14_out=8'h3e;
		8'h6d: mul14_out=8'h30;
		8'h6e: mul14_out=8'h22;
		8'h6f: mul14_out=8'h2c;
		8'h70: mul14_out=8'h96;
		8'h71: mul14_out=8'h98;
		8'h72: mul14_out=8'h8a;
		8'h73: mul14_out=8'h84;
		8'h74: mul14_out=8'hae;
		8'h75: mul14_out=8'ha0;
		8'h76: mul14_out=8'hb2;
		8'h77: mul14_out=8'hbc;
		8'h78: mul14_out=8'he6;
		8'h79: mul14_out=8'he8;
		8'h7a: mul14_out=8'hfa;
		8'h7b: mul14_out=8'hf4;
		8'h7c: mul14_out=8'hde;
		8'h7d: mul14_out=8'hd0;
		8'h7e: mul14_out=8'hc2;
		8'h7f: mul14_out=8'hcc;
		8'h80: mul14_out=8'h41;
		8'h81: mul14_out=8'h4f;
		8'h82: mul14_out=8'h5d;
		8'h83: mul14_out=8'h53;
		8'h84: mul14_out=8'h79;
		8'h85: mul14_out=8'h77;
		8'h86: mul14_out=8'h65;
		8'h87: mul14_out=8'h6b;
		8'h88: mul14_out=8'h31;
		8'h89: mul14_out=8'h3f;
		8'h8a: mul14_out=8'h2d;
		8'h8b: mul14_out=8'h23;
		8'h8c: mul14_out=8'h09;
		8'h8d: mul14_out=8'h07;
		8'h8e: mul14_out=8'h15;
		8'h8f: mul14_out=8'h1b;
		8'h90: mul14_out=8'ha1;
		8'h91: mul14_out=8'haf;
		8'h92: mul14_out=8'hbd;
		8'h93: mul14_out=8'hb3;
		8'h94: mul14_out=8'h99;
		8'h95: mul14_out=8'h97;
		8'h96: mul14_out=8'h85;
		8'h97: mul14_out=8'h8b;
		8'h98: mul14_out=8'hd1;
		8'h99: mul14_out=8'hdf;
		8'h9a: mul14_out=8'hcd;
		8'h9b: mul14_out=8'hc3;
		8'h9c: mul14_out=8'he9;
		8'h9d: mul14_out=8'he7;
		8'h9e: mul14_out=8'hf5;
		8'h9f: mul14_out=8'hfb;
		8'ha0: mul14_out=8'h9a;
		8'ha1: mul14_out=8'h94;
		8'ha2: mul14_out=8'h86;
		8'ha3: mul14_out=8'h88;
		8'ha4: mul14_out=8'ha2;
		8'ha5: mul14_out=8'hac;
		8'ha6: mul14_out=8'hbe;
		8'ha7: mul14_out=8'hb0;
		8'ha8: mul14_out=8'hea;
		8'ha9: mul14_out=8'he4;
		8'haa: mul14_out=8'hf6;
		8'hab: mul14_out=8'hf8;
		8'hac: mul14_out=8'hd2;
		8'had: mul14_out=8'hdc;
		8'hae: mul14_out=8'hce;
		8'haf: mul14_out=8'hc0;
		8'hb0: mul14_out=8'h7a;
		8'hb1: mul14_out=8'h74;
		8'hb2: mul14_out=8'h66;
		8'hb3: mul14_out=8'h68;
		8'hb4: mul14_out=8'h42;
		8'hb5: mul14_out=8'h4c;
		8'hb6: mul14_out=8'h5e;
		8'hb7: mul14_out=8'h50;
		8'hb8: mul14_out=8'h0a;
		8'hb9: mul14_out=8'h04;
		8'hba: mul14_out=8'h16;
		8'hbb: mul14_out=8'h18;
		8'hbc: mul14_out=8'h32;
		8'hbd: mul14_out=8'h3c;
		8'hbe: mul14_out=8'h2e;
		8'hbf: mul14_out=8'h20;
		8'hc0: mul14_out=8'hec;
		8'hc1: mul14_out=8'he2;
		8'hc2: mul14_out=8'hf0;
		8'hc3: mul14_out=8'hfe;
		8'hc4: mul14_out=8'hd4;
		8'hc5: mul14_out=8'hda;
		8'hc6: mul14_out=8'hc8;
		8'hc7: mul14_out=8'hc6;
		8'hc8: mul14_out=8'h9c;
		8'hc9: mul14_out=8'h92;
		8'hca: mul14_out=8'h80;
		8'hcb: mul14_out=8'h8e;
		8'hcc: mul14_out=8'ha4;
		8'hcd: mul14_out=8'haa;
		8'hce: mul14_out=8'hb8;
		8'hcf: mul14_out=8'hb6;
		8'hd0: mul14_out=8'h0c;
		8'hd1: mul14_out=8'h02;
		8'hd2: mul14_out=8'h10;
		8'hd3: mul14_out=8'h1e;
		8'hd4: mul14_out=8'h34;
		8'hd5: mul14_out=8'h3a;
		8'hd6: mul14_out=8'h28;
		8'hd7: mul14_out=8'h26;
		8'hd8: mul14_out=8'h7c;
		8'hd9: mul14_out=8'h72;
		8'hda: mul14_out=8'h60;
		8'hdb: mul14_out=8'h6e;
		8'hdc: mul14_out=8'h44;
		8'hdd: mul14_out=8'h4a;
		8'hde: mul14_out=8'h58;
		8'hdf: mul14_out=8'h56;
		8'he0: mul14_out=8'h37;
		8'he1: mul14_out=8'h39;
		8'he2: mul14_out=8'h2b;
		8'he3: mul14_out=8'h25;
		8'he4: mul14_out=8'h0f;
		8'he5: mul14_out=8'h01;
		8'he6: mul14_out=8'h13;
		8'he7: mul14_out=8'h1d;
		8'he8: mul14_out=8'h47;
		8'he9: mul14_out=8'h49;
		8'hea: mul14_out=8'h5b;
		8'heb: mul14_out=8'h55;
		8'hec: mul14_out=8'h7f;
		8'hed: mul14_out=8'h71;
		8'hee: mul14_out=8'h63;
		8'hef: mul14_out=8'h6d;
		8'hf0: mul14_out=8'hd7;
		8'hf1: mul14_out=8'hd9;
		8'hf2: mul14_out=8'hcb;
		8'hf3: mul14_out=8'hc5;
		8'hf4: mul14_out=8'hef;
		8'hf5: mul14_out=8'he1;
		8'hf6: mul14_out=8'hf3;
		8'hf7: mul14_out=8'hfd;
		8'hf8: mul14_out=8'ha7;
		8'hf9: mul14_out=8'ha9;
		8'hfa: mul14_out=8'hbb;
		8'hfb: mul14_out=8'hb5;
		8'hfc: mul14_out=8'h9f;
		8'hfd: mul14_out=8'h91;
		8'hfe: mul14_out=8'h83;
		8'hff: mul14_out=8'h8d;
endcase
end

endmodule
