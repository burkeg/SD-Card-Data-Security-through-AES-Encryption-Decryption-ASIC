// $Id: $
// File name:   i_s_box.sv
// Created:     3/12/2017
// Author:      Gabriel Burke
// Lab Section: 337-02
// Version:     1.0  Initial Design Entry
// Description: Inverse Rijndael S-Box 

module i_s_box(
	input wire [7:0]i_s_box_in,
	output reg [7:0]i_s_box_out
);

always_comb begin : i_s_box_case
	i_s_box_out=8'h63;

	case(i_s_box_in)
	8'h00: i_s_box_out=8'h52;
	8'h01: i_s_box_out=8'h09;
	8'h02: i_s_box_out=8'h6a;
	8'h03: i_s_box_out=8'hd5;
	8'h04: i_s_box_out=8'h30;
	8'h05: i_s_box_out=8'h36;
	8'h06: i_s_box_out=8'ha5;
	8'h07: i_s_box_out=8'h38;
	8'h08: i_s_box_out=8'hbf;
	8'h09: i_s_box_out=8'h40;
	8'h0a: i_s_box_out=8'ha3;
	8'h0b: i_s_box_out=8'h9e;
	8'h0c: i_s_box_out=8'h81;
	8'h0d: i_s_box_out=8'hf3;
	8'h0e: i_s_box_out=8'hd7;
	8'h0f: i_s_box_out=8'hfb;
	8'h10: i_s_box_out=8'h7c;
	8'h11: i_s_box_out=8'he3;
	8'h12: i_s_box_out=8'h39;
	8'h13: i_s_box_out=8'h82;
	8'h14: i_s_box_out=8'h9b;
	8'h15: i_s_box_out=8'h2f;
	8'h16: i_s_box_out=8'hff;
	8'h17: i_s_box_out=8'h87;
	8'h18: i_s_box_out=8'h34;
	8'h19: i_s_box_out=8'h8e;
	8'h1a: i_s_box_out=8'h43;
	8'h1b: i_s_box_out=8'h44;
	8'h1c: i_s_box_out=8'hc4;
	8'h1d: i_s_box_out=8'hde;
	8'h1e: i_s_box_out=8'he9;
	8'h1f: i_s_box_out=8'hcb;
	8'h20: i_s_box_out=8'h54;
	8'h21: i_s_box_out=8'h7b;
	8'h22: i_s_box_out=8'h94;
	8'h23: i_s_box_out=8'h32;
	8'h24: i_s_box_out=8'ha6;
	8'h25: i_s_box_out=8'hc2;
	8'h26: i_s_box_out=8'h23;
	8'h27: i_s_box_out=8'h3d;
	8'h28: i_s_box_out=8'hee;
	8'h29: i_s_box_out=8'h4c;
	8'h2a: i_s_box_out=8'h95;
	8'h2b: i_s_box_out=8'h0b;
	8'h2c: i_s_box_out=8'h42;
	8'h2d: i_s_box_out=8'hfa;
	8'h2e: i_s_box_out=8'hc3;
	8'h2f: i_s_box_out=8'h4e;
	8'h30: i_s_box_out=8'h08;
	8'h31: i_s_box_out=8'h2e;
	8'h32: i_s_box_out=8'ha1;
	8'h33: i_s_box_out=8'h66;
	8'h34: i_s_box_out=8'h28;
	8'h35: i_s_box_out=8'hd9;
	8'h36: i_s_box_out=8'h24;
	8'h37: i_s_box_out=8'hb2;
	8'h38: i_s_box_out=8'h76;
	8'h39: i_s_box_out=8'h5b;
	8'h3a: i_s_box_out=8'ha2;
	8'h3b: i_s_box_out=8'h49;
	8'h3c: i_s_box_out=8'h6d;
	8'h3d: i_s_box_out=8'h8b;
	8'h3e: i_s_box_out=8'hd1;
	8'h3f: i_s_box_out=8'h25;
	8'h40: i_s_box_out=8'h72;
	8'h41: i_s_box_out=8'hf8;
	8'h42: i_s_box_out=8'hf6;
	8'h43: i_s_box_out=8'h64;
	8'h44: i_s_box_out=8'h86;
	8'h45: i_s_box_out=8'h68;
	8'h46: i_s_box_out=8'h98;
	8'h47: i_s_box_out=8'h16;
	8'h48: i_s_box_out=8'hd4;
	8'h49: i_s_box_out=8'ha4;
	8'h4a: i_s_box_out=8'h5c;
	8'h4b: i_s_box_out=8'hcc;
	8'h4c: i_s_box_out=8'h5d;
	8'h4d: i_s_box_out=8'h65;
	8'h4e: i_s_box_out=8'hb6;
	8'h4f: i_s_box_out=8'h92;
	8'h50: i_s_box_out=8'h6c;
	8'h51: i_s_box_out=8'h70;
	8'h52: i_s_box_out=8'h48;
	8'h53: i_s_box_out=8'h50;
	8'h54: i_s_box_out=8'hfd;
	8'h55: i_s_box_out=8'hed;
	8'h56: i_s_box_out=8'hb9;
	8'h57: i_s_box_out=8'hda;
	8'h58: i_s_box_out=8'h5e;
	8'h59: i_s_box_out=8'h15;
	8'h5a: i_s_box_out=8'h46;
	8'h5b: i_s_box_out=8'h57;
	8'h5c: i_s_box_out=8'ha7;
	8'h5d: i_s_box_out=8'h8d;
	8'h5e: i_s_box_out=8'h9d;
	8'h5f: i_s_box_out=8'h84;
	8'h60: i_s_box_out=8'h90;
	8'h61: i_s_box_out=8'hd8;
	8'h62: i_s_box_out=8'hab;
	8'h63: i_s_box_out=8'h00;
	8'h64: i_s_box_out=8'h8c;
	8'h65: i_s_box_out=8'hbc;
	8'h66: i_s_box_out=8'hd3;
	8'h67: i_s_box_out=8'h0a;
	8'h68: i_s_box_out=8'hf7;
	8'h69: i_s_box_out=8'he4;
	8'h6a: i_s_box_out=8'h58;
	8'h6b: i_s_box_out=8'h05;
	8'h6c: i_s_box_out=8'hb8;
	8'h6d: i_s_box_out=8'hb3;
	8'h6e: i_s_box_out=8'h45;
	8'h6f: i_s_box_out=8'h06;
	8'h70: i_s_box_out=8'hd0;
	8'h71: i_s_box_out=8'h2c;
	8'h72: i_s_box_out=8'h1e;
	8'h73: i_s_box_out=8'h8f;
	8'h74: i_s_box_out=8'hca;
	8'h75: i_s_box_out=8'h3f;
	8'h76: i_s_box_out=8'h0f;
	8'h77: i_s_box_out=8'h02;
	8'h78: i_s_box_out=8'hc1;
	8'h79: i_s_box_out=8'haf;
	8'h7a: i_s_box_out=8'hbd;
	8'h7b: i_s_box_out=8'h03;
	8'h7c: i_s_box_out=8'h01;
	8'h7d: i_s_box_out=8'h13;
	8'h7e: i_s_box_out=8'h8a;
	8'h7f: i_s_box_out=8'h6b;
	8'h80: i_s_box_out=8'h3a;
	8'h81: i_s_box_out=8'h91;
	8'h82: i_s_box_out=8'h11;
	8'h83: i_s_box_out=8'h41;
	8'h84: i_s_box_out=8'h4f;
	8'h85: i_s_box_out=8'h67;
	8'h86: i_s_box_out=8'hdc;
	8'h87: i_s_box_out=8'hea;
	8'h88: i_s_box_out=8'h97;
	8'h89: i_s_box_out=8'hf2;
	8'h8a: i_s_box_out=8'hcf;
	8'h8b: i_s_box_out=8'hce;
	8'h8c: i_s_box_out=8'hf0;
	8'h8d: i_s_box_out=8'hb4;
	8'h8e: i_s_box_out=8'he6;
	8'h8f: i_s_box_out=8'h73;
	8'h90: i_s_box_out=8'h96;
	8'h91: i_s_box_out=8'hac;
	8'h92: i_s_box_out=8'h74;
	8'h93: i_s_box_out=8'h22;
	8'h94: i_s_box_out=8'he7;
	8'h95: i_s_box_out=8'had;
	8'h96: i_s_box_out=8'h35;
	8'h97: i_s_box_out=8'h85;
	8'h98: i_s_box_out=8'he2;
	8'h99: i_s_box_out=8'hf9;
	8'h9a: i_s_box_out=8'h37;
	8'h9b: i_s_box_out=8'he8;
	8'h9c: i_s_box_out=8'h1c;
	8'h9d: i_s_box_out=8'h75;
	8'h9e: i_s_box_out=8'hdf;
	8'h9f: i_s_box_out=8'h6e;
	8'ha0: i_s_box_out=8'h47;
	8'ha1: i_s_box_out=8'hf1;
	8'ha2: i_s_box_out=8'h1a;
	8'ha3: i_s_box_out=8'h71;
	8'ha4: i_s_box_out=8'h1d;
	8'ha5: i_s_box_out=8'h29;
	8'ha6: i_s_box_out=8'hc5;
	8'ha7: i_s_box_out=8'h89;
	8'ha8: i_s_box_out=8'h6f;
	8'ha9: i_s_box_out=8'hb7;
	8'haa: i_s_box_out=8'h62;
	8'hab: i_s_box_out=8'h0e;
	8'hac: i_s_box_out=8'haa;
	8'had: i_s_box_out=8'h18;
	8'hae: i_s_box_out=8'hbe;
	8'haf: i_s_box_out=8'h1b;
	8'hb0: i_s_box_out=8'hfc;
	8'hb1: i_s_box_out=8'h56;
	8'hb2: i_s_box_out=8'h3e;
	8'hb3: i_s_box_out=8'h4b;
	8'hb4: i_s_box_out=8'hc6;
	8'hb5: i_s_box_out=8'hd2;
	8'hb6: i_s_box_out=8'h79;
	8'hb7: i_s_box_out=8'h20;
	8'hb8: i_s_box_out=8'h9a;
	8'hb9: i_s_box_out=8'hdb;
	8'hba: i_s_box_out=8'hc0;
	8'hbb: i_s_box_out=8'hfe;
	8'hbc: i_s_box_out=8'h78;
	8'hbd: i_s_box_out=8'hcd;
	8'hbe: i_s_box_out=8'h5a;
	8'hbf: i_s_box_out=8'hf4;
	8'hc0: i_s_box_out=8'h1f;
	8'hc1: i_s_box_out=8'hdd;
	8'hc2: i_s_box_out=8'ha8;
	8'hc3: i_s_box_out=8'h33;
	8'hc4: i_s_box_out=8'h88;
	8'hc5: i_s_box_out=8'h07;
	8'hc6: i_s_box_out=8'hc7;
	8'hc7: i_s_box_out=8'h31;
	8'hc8: i_s_box_out=8'hb1;
	8'hc9: i_s_box_out=8'h12;
	8'hca: i_s_box_out=8'h10;
	8'hcb: i_s_box_out=8'h59;
	8'hcc: i_s_box_out=8'h27;
	8'hcd: i_s_box_out=8'h80;
	8'hce: i_s_box_out=8'hec;
	8'hcf: i_s_box_out=8'h5f;
	8'hd0: i_s_box_out=8'h60;
	8'hd1: i_s_box_out=8'h51;
	8'hd2: i_s_box_out=8'h7f;
	8'hd3: i_s_box_out=8'ha9;
	8'hd4: i_s_box_out=8'h19;
	8'hd5: i_s_box_out=8'hb5;
	8'hd6: i_s_box_out=8'h4a;
	8'hd7: i_s_box_out=8'h0d;
	8'hd8: i_s_box_out=8'h2d;
	8'hd9: i_s_box_out=8'he5;
	8'hda: i_s_box_out=8'h7a;
	8'hdb: i_s_box_out=8'h9f;
	8'hdc: i_s_box_out=8'h93;
	8'hdd: i_s_box_out=8'hc9;
	8'hde: i_s_box_out=8'h9c;
	8'hdf: i_s_box_out=8'hef;
	8'he0: i_s_box_out=8'ha0;
	8'he1: i_s_box_out=8'he0;
	8'he2: i_s_box_out=8'h3b;
	8'he3: i_s_box_out=8'h4d;
	8'he4: i_s_box_out=8'hae;
	8'he5: i_s_box_out=8'h2a;
	8'he6: i_s_box_out=8'hf5;
	8'he7: i_s_box_out=8'hb0;
	8'he8: i_s_box_out=8'hc8;
	8'he9: i_s_box_out=8'heb;
	8'hea: i_s_box_out=8'hbb;
	8'heb: i_s_box_out=8'h3c;
	8'hec: i_s_box_out=8'h83;
	8'hed: i_s_box_out=8'h53;
	8'hee: i_s_box_out=8'h99;
	8'hef: i_s_box_out=8'h61;
	8'hf0: i_s_box_out=8'h17;
	8'hf1: i_s_box_out=8'h2b;
	8'hf2: i_s_box_out=8'h04;
	8'hf3: i_s_box_out=8'h7e;
	8'hf4: i_s_box_out=8'hba;
	8'hf5: i_s_box_out=8'h77;
	8'hf6: i_s_box_out=8'hd6;
	8'hf7: i_s_box_out=8'h26;
	8'hf8: i_s_box_out=8'he1;
	8'hf9: i_s_box_out=8'h69;
	8'hfa: i_s_box_out=8'h14;
	8'hfb: i_s_box_out=8'h63;
	8'hfc: i_s_box_out=8'h55;
	8'hfd: i_s_box_out=8'h21;
	8'hfe: i_s_box_out=8'h0c;
	8'hff: i_s_box_out=8'h7d;
endcase
end

endmodule